// pfl_fl.v

// Generated using ACDS version 14.0 200 at 2015.07.15.09:35:40

`timescale 1 ps / 1 ps
module pfl_fl (
		input  wire        pfl_nreset,               //               pfl_nreset.pfl_nreset
		input  wire        pfl_flash_access_granted, // pfl_flash_access_granted.pfl_flash_access_granted
		output wire        pfl_flash_access_request, // pfl_flash_access_request.pfl_flash_access_request
		output wire [24:0] flash_addr,               //               flash_addr.flash_addr
		inout  wire [15:0] flash_data,               //               flash_data.flash_data
		output wire        flash_nce,                //                flash_nce.flash_nce
		output wire        flash_nwe,                //                flash_nwe.flash_nwe
		output wire        flash_noe,                //                flash_noe.flash_noe
		input  wire        pfl_clk,                  //                  pfl_clk.pfl_clk
		input  wire [2:0]  fpga_pgm,                 //                 fpga_pgm.fpga_pgm
		input  wire        fpga_conf_done,           //           fpga_conf_done.fpga_conf_done
		input  wire        fpga_nstatus,             //             fpga_nstatus.fpga_nstatus
		output wire        fpga_data,                //                fpga_data.fpga_data
		output wire        fpga_dclk,                //                fpga_dclk.fpga_dclk
		output wire        fpga_nconfig              //             fpga_nconfig.fpga_nconfig
	);

	altera_parallel_flash_loader #(
		.TRISTATE_CHECKBOX          (1),
		.FEATURES_PGM               (1),
		.FEATURES_CFG               (1),
		.FLASH_TYPE                 ("CFI_FLASH"),
		.ADDR_WIDTH                 (25),
		.FLASH_DATA_WIDTH           (16),
		.N_FLASH                    (1),
		.FLASH_NRESET_CHECKBOX      (0),
		.ENHANCED_FLASH_PROGRAMMING (0),
		.FIFO_SIZE                  (16),
		.DISABLE_CRC_CHECKBOX       (0),
		.CLK_DIVISOR                (9),
		.PAGE_CLK_DIVISOR           (2),
		.FLASH_NRESET_COUNTER       (5000),
		.NORMAL_MODE                (1),
		.BURST_MODE                 (0),
		.PAGE_MODE                  (0),
		.BURST_MODE_SPANSION        (0),
		.BURST_MODE_INTEL           (0),
		.BURST_MODE_LATENCY_COUNT   (3),
		.BURST_MODE_NUMONYX         (0),
		.FLASH_BURST_EXTRA_CYCLE    (1),
		.CONF_DATA_WIDTH            (1),
		.OPTION_BITS_START_ADDRESS  (0),
		.CONF_WAIT_TIMER_WIDTH      (20),
		.DCLK_DIVISOR               (1),
		.DECOMPRESSOR_MODE          ("NONE"),
		.SAFE_MODE_HALT             (1),
		.SAFE_MODE_RETRY            (0),
		.SAFE_MODE_REVERT           (0),
		.SAFE_MODE_REVERT_ADDR      (0),
		.QSPI_DATA_DELAY            (0),
		.QSPI_DATA_DELAY_COUNT      (1)
	) parallel_flash_loader_0 (
		.pfl_nreset               (pfl_nreset),               //               pfl_nreset.pfl_nreset
		.pfl_flash_access_granted (pfl_flash_access_granted), // pfl_flash_access_granted.pfl_flash_access_granted
		.pfl_clk                  (pfl_clk),                  //                  pfl_clk.pfl_clk
		.fpga_pgm                 (fpga_pgm),                 //                 fpga_pgm.fpga_pgm
		.fpga_conf_done           (fpga_conf_done),           //           fpga_conf_done.fpga_conf_done
		.fpga_nstatus             (fpga_nstatus),             //             fpga_nstatus.fpga_nstatus
		.pfl_flash_access_request (pfl_flash_access_request), // pfl_flash_access_request.pfl_flash_access_request
		.flash_addr               (flash_addr),               //               flash_addr.flash_addr
		.flash_data               (flash_data),               //               flash_data.flash_data
		.flash_nce                (flash_nce),                //                flash_nce.flash_nce
		.flash_nwe                (flash_nwe),                //                flash_nwe.flash_nwe
		.flash_noe                (flash_noe),                //                flash_noe.flash_noe
		.fpga_data                (fpga_data),                //                fpga_data.fpga_data
		.fpga_dclk                (fpga_dclk),                //                fpga_dclk.fpga_dclk
		.fpga_nconfig             (fpga_nconfig)              //             fpga_nconfig.fpga_nconfig
	);

endmodule
